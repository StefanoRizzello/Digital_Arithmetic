federica@federica-X556URK.18911:1637582398